module sll(data_operandA, ctrl_shiftamt, shifted_output, shift_enable);

	input [31:0] data_operandA;
	input [4:0] ctrl_shiftamt;
	input shift_enable;
	wire [31:0] muxed_output;
	output [31:0] shifted_output;
	
	wire [31:0] in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31;
	
	mux_32 mux_32_sll(muxed_output, ctrl_shiftamt, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31);
	
	and and_0(shifted_output[0], muxed_output[0], shift_enable);
	and and_1(shifted_output[1], muxed_output[1], shift_enable);
	and and_2(shifted_output[2], muxed_output[2], shift_enable);
	and and_3(shifted_output[3], muxed_output[3], shift_enable);
	and and_4(shifted_output[4], muxed_output[4], shift_enable);
	and and_5(shifted_output[5], muxed_output[5], shift_enable);
	and and_6(shifted_output[6], muxed_output[6], shift_enable);
	and and_7(shifted_output[7], muxed_output[7], shift_enable);
	and and_8(shifted_output[8], muxed_output[8], shift_enable);
	and and_9(shifted_output[9], muxed_output[9], shift_enable);
	and and_10(shifted_output[10], muxed_output[10], shift_enable);
	and and_11(shifted_output[11], muxed_output[11], shift_enable);
	and and_12(shifted_output[12], muxed_output[12], shift_enable);
	and and_13(shifted_output[13], muxed_output[13], shift_enable);
	and and_14(shifted_output[14], muxed_output[14], shift_enable);
	and and_15(shifted_output[15], muxed_output[15], shift_enable);
	and and_16(shifted_output[16], muxed_output[16], shift_enable);
	and and_17(shifted_output[17], muxed_output[17], shift_enable);
	and and_18(shifted_output[18], muxed_output[18], shift_enable);
	and and_19(shifted_output[19], muxed_output[19], shift_enable);
	and and_20(shifted_output[20], muxed_output[20], shift_enable);
	and and_21(shifted_output[21], muxed_output[21], shift_enable);
	and and_22(shifted_output[22], muxed_output[22], shift_enable);
	and and_23(shifted_output[23], muxed_output[23], shift_enable);
	and and_24(shifted_output[24], muxed_output[24], shift_enable);
	and and_25(shifted_output[25], muxed_output[25], shift_enable);
	and and_26(shifted_output[26], muxed_output[26], shift_enable);
	and and_27(shifted_output[27], muxed_output[27], shift_enable);
	and and_28(shifted_output[28], muxed_output[28], shift_enable);
	and and_29(shifted_output[29], muxed_output[29], shift_enable);
	and and_30(shifted_output[30], muxed_output[30], shift_enable);
	and and_31(shifted_output[31], muxed_output[31], shift_enable);
	
assign in0[31:0] = data_operandA[31:0];
assign in1[31:1] = data_operandA[30:0];
assign in1[0] = 0;
assign in2[31:2] = data_operandA[29:0];
assign in2[0] = 0;
assign in2[1] = 0;
assign in3[31:3] = data_operandA[28:0];
assign in3[0] = 0;
assign in3[1] = 0;
assign in3[2] = 0;
assign in4[31:4] = data_operandA[27:0];
assign in4[0] = 0;
assign in4[1] = 0;
assign in4[2] = 0;
assign in4[3] = 0;
assign in5[31:5] = data_operandA[26:0];
assign in5[0] = 0;
assign in5[1] = 0;
assign in5[2] = 0;
assign in5[3] = 0;
assign in5[4] = 0;
assign in6[31:6] = data_operandA[25:0];
assign in6[0] = 0;
assign in6[1] = 0;
assign in6[2] = 0;
assign in6[3] = 0;
assign in6[4] = 0;
assign in6[5] = 0;
assign in7[31:7] = data_operandA[24:0];
assign in7[0] = 0;
assign in7[1] = 0;
assign in7[2] = 0;
assign in7[3] = 0;
assign in7[4] = 0;
assign in7[5] = 0;
assign in7[6] = 0;
assign in8[31:8] = data_operandA[23:0];
assign in8[0] = 0;
assign in8[1] = 0;
assign in8[2] = 0;
assign in8[3] = 0;
assign in8[4] = 0;
assign in8[5] = 0;
assign in8[6] = 0;
assign in8[7] = 0;
assign in9[31:9] = data_operandA[22:0];
assign in9[0] = 0;
assign in9[1] = 0;
assign in9[2] = 0;
assign in9[3] = 0;
assign in9[4] = 0;
assign in9[5] = 0;
assign in9[6] = 0;
assign in9[7] = 0;
assign in9[8] = 0;
assign in10[31:10] = data_operandA[21:0];
assign in10[0] = 0;
assign in10[1] = 0;
assign in10[2] = 0;
assign in10[3] = 0;
assign in10[4] = 0;
assign in10[5] = 0;
assign in10[6] = 0;
assign in10[7] = 0;
assign in10[8] = 0;
assign in10[9] = 0;
assign in11[31:11] = data_operandA[20:0];
assign in11[0] = 0;
assign in11[1] = 0;
assign in11[2] = 0;
assign in11[3] = 0;
assign in11[4] = 0;
assign in11[5] = 0;
assign in11[6] = 0;
assign in11[7] = 0;
assign in11[8] = 0;
assign in11[9] = 0;
assign in11[10] = 0;
assign in12[31:12] = data_operandA[19:0];
assign in12[0] = 0;
assign in12[1] = 0;
assign in12[2] = 0;
assign in12[3] = 0;
assign in12[4] = 0;
assign in12[5] = 0;
assign in12[6] = 0;
assign in12[7] = 0;
assign in12[8] = 0;
assign in12[9] = 0;
assign in12[10] = 0;
assign in12[11] = 0;
assign in13[31:13] = data_operandA[18:0];
assign in13[0] = 0;
assign in13[1] = 0;
assign in13[2] = 0;
assign in13[3] = 0;
assign in13[4] = 0;
assign in13[5] = 0;
assign in13[6] = 0;
assign in13[7] = 0;
assign in13[8] = 0;
assign in13[9] = 0;
assign in13[10] = 0;
assign in13[11] = 0;
assign in13[12] = 0;
assign in14[31:14] = data_operandA[17:0];
assign in14[0] = 0;
assign in14[1] = 0;
assign in14[2] = 0;
assign in14[3] = 0;
assign in14[4] = 0;
assign in14[5] = 0;
assign in14[6] = 0;
assign in14[7] = 0;
assign in14[8] = 0;
assign in14[9] = 0;
assign in14[10] = 0;
assign in14[11] = 0;
assign in14[12] = 0;
assign in14[13] = 0;
assign in15[31:15] = data_operandA[16:0];
assign in15[0] = 0;
assign in15[1] = 0;
assign in15[2] = 0;
assign in15[3] = 0;
assign in15[4] = 0;
assign in15[5] = 0;
assign in15[6] = 0;
assign in15[7] = 0;
assign in15[8] = 0;
assign in15[9] = 0;
assign in15[10] = 0;
assign in15[11] = 0;
assign in15[12] = 0;
assign in15[13] = 0;
assign in15[14] = 0;
assign in16[31:16] = data_operandA[15:0];
assign in16[0] = 0;
assign in16[1] = 0;
assign in16[2] = 0;
assign in16[3] = 0;
assign in16[4] = 0;
assign in16[5] = 0;
assign in16[6] = 0;
assign in16[7] = 0;
assign in16[8] = 0;
assign in16[9] = 0;
assign in16[10] = 0;
assign in16[11] = 0;
assign in16[12] = 0;
assign in16[13] = 0;
assign in16[14] = 0;
assign in16[15] = 0;
assign in17[31:17] = data_operandA[14:0];
assign in17[0] = 0;
assign in17[1] = 0;
assign in17[2] = 0;
assign in17[3] = 0;
assign in17[4] = 0;
assign in17[5] = 0;
assign in17[6] = 0;
assign in17[7] = 0;
assign in17[8] = 0;
assign in17[9] = 0;
assign in17[10] = 0;
assign in17[11] = 0;
assign in17[12] = 0;
assign in17[13] = 0;
assign in17[14] = 0;
assign in17[15] = 0;
assign in17[16] = 0;
assign in18[31:18] = data_operandA[13:0];
assign in18[0] = 0;
assign in18[1] = 0;
assign in18[2] = 0;
assign in18[3] = 0;
assign in18[4] = 0;
assign in18[5] = 0;
assign in18[6] = 0;
assign in18[7] = 0;
assign in18[8] = 0;
assign in18[9] = 0;
assign in18[10] = 0;
assign in18[11] = 0;
assign in18[12] = 0;
assign in18[13] = 0;
assign in18[14] = 0;
assign in18[15] = 0;
assign in18[16] = 0;
assign in18[17] = 0;
assign in19[31:19] = data_operandA[12:0];
assign in19[0] = 0;
assign in19[1] = 0;
assign in19[2] = 0;
assign in19[3] = 0;
assign in19[4] = 0;
assign in19[5] = 0;
assign in19[6] = 0;
assign in19[7] = 0;
assign in19[8] = 0;
assign in19[9] = 0;
assign in19[10] = 0;
assign in19[11] = 0;
assign in19[12] = 0;
assign in19[13] = 0;
assign in19[14] = 0;
assign in19[15] = 0;
assign in19[16] = 0;
assign in19[17] = 0;
assign in19[18] = 0;
assign in20[31:20] = data_operandA[11:0];
assign in20[0] = 0;
assign in20[1] = 0;
assign in20[2] = 0;
assign in20[3] = 0;
assign in20[4] = 0;
assign in20[5] = 0;
assign in20[6] = 0;
assign in20[7] = 0;
assign in20[8] = 0;
assign in20[9] = 0;
assign in20[10] = 0;
assign in20[11] = 0;
assign in20[12] = 0;
assign in20[13] = 0;
assign in20[14] = 0;
assign in20[15] = 0;
assign in20[16] = 0;
assign in20[17] = 0;
assign in20[18] = 0;
assign in20[19] = 0;
assign in21[31:21] = data_operandA[10:0];
assign in21[0] = 0;
assign in21[1] = 0;
assign in21[2] = 0;
assign in21[3] = 0;
assign in21[4] = 0;
assign in21[5] = 0;
assign in21[6] = 0;
assign in21[7] = 0;
assign in21[8] = 0;
assign in21[9] = 0;
assign in21[10] = 0;
assign in21[11] = 0;
assign in21[12] = 0;
assign in21[13] = 0;
assign in21[14] = 0;
assign in21[15] = 0;
assign in21[16] = 0;
assign in21[17] = 0;
assign in21[18] = 0;
assign in21[19] = 0;
assign in21[20] = 0;
assign in22[31:22] = data_operandA[9:0];
assign in22[0] = 0;
assign in22[1] = 0;
assign in22[2] = 0;
assign in22[3] = 0;
assign in22[4] = 0;
assign in22[5] = 0;
assign in22[6] = 0;
assign in22[7] = 0;
assign in22[8] = 0;
assign in22[9] = 0;
assign in22[10] = 0;
assign in22[11] = 0;
assign in22[12] = 0;
assign in22[13] = 0;
assign in22[14] = 0;
assign in22[15] = 0;
assign in22[16] = 0;
assign in22[17] = 0;
assign in22[18] = 0;
assign in22[19] = 0;
assign in22[20] = 0;
assign in22[21] = 0;
assign in23[31:23] = data_operandA[8:0];
assign in23[0] = 0;
assign in23[1] = 0;
assign in23[2] = 0;
assign in23[3] = 0;
assign in23[4] = 0;
assign in23[5] = 0;
assign in23[6] = 0;
assign in23[7] = 0;
assign in23[8] = 0;
assign in23[9] = 0;
assign in23[10] = 0;
assign in23[11] = 0;
assign in23[12] = 0;
assign in23[13] = 0;
assign in23[14] = 0;
assign in23[15] = 0;
assign in23[16] = 0;
assign in23[17] = 0;
assign in23[18] = 0;
assign in23[19] = 0;
assign in23[20] = 0;
assign in23[21] = 0;
assign in23[22] = 0;
assign in24[31:24] = data_operandA[7:0];
assign in24[0] = 0;
assign in24[1] = 0;
assign in24[2] = 0;
assign in24[3] = 0;
assign in24[4] = 0;
assign in24[5] = 0;
assign in24[6] = 0;
assign in24[7] = 0;
assign in24[8] = 0;
assign in24[9] = 0;
assign in24[10] = 0;
assign in24[11] = 0;
assign in24[12] = 0;
assign in24[13] = 0;
assign in24[14] = 0;
assign in24[15] = 0;
assign in24[16] = 0;
assign in24[17] = 0;
assign in24[18] = 0;
assign in24[19] = 0;
assign in24[20] = 0;
assign in24[21] = 0;
assign in24[22] = 0;
assign in24[23] = 0;
assign in25[31:25] = data_operandA[6:0];
assign in25[0] = 0;
assign in25[1] = 0;
assign in25[2] = 0;
assign in25[3] = 0;
assign in25[4] = 0;
assign in25[5] = 0;
assign in25[6] = 0;
assign in25[7] = 0;
assign in25[8] = 0;
assign in25[9] = 0;
assign in25[10] = 0;
assign in25[11] = 0;
assign in25[12] = 0;
assign in25[13] = 0;
assign in25[14] = 0;
assign in25[15] = 0;
assign in25[16] = 0;
assign in25[17] = 0;
assign in25[18] = 0;
assign in25[19] = 0;
assign in25[20] = 0;
assign in25[21] = 0;
assign in25[22] = 0;
assign in25[23] = 0;
assign in25[24] = 0;
assign in26[31:26] = data_operandA[5:0];
assign in26[0] = 0;
assign in26[1] = 0;
assign in26[2] = 0;
assign in26[3] = 0;
assign in26[4] = 0;
assign in26[5] = 0;
assign in26[6] = 0;
assign in26[7] = 0;
assign in26[8] = 0;
assign in26[9] = 0;
assign in26[10] = 0;
assign in26[11] = 0;
assign in26[12] = 0;
assign in26[13] = 0;
assign in26[14] = 0;
assign in26[15] = 0;
assign in26[16] = 0;
assign in26[17] = 0;
assign in26[18] = 0;
assign in26[19] = 0;
assign in26[20] = 0;
assign in26[21] = 0;
assign in26[22] = 0;
assign in26[23] = 0;
assign in26[24] = 0;
assign in26[25] = 0;
assign in27[31:27] = data_operandA[4:0];
assign in27[0] = 0;
assign in27[1] = 0;
assign in27[2] = 0;
assign in27[3] = 0;
assign in27[4] = 0;
assign in27[5] = 0;
assign in27[6] = 0;
assign in27[7] = 0;
assign in27[8] = 0;
assign in27[9] = 0;
assign in27[10] = 0;
assign in27[11] = 0;
assign in27[12] = 0;
assign in27[13] = 0;
assign in27[14] = 0;
assign in27[15] = 0;
assign in27[16] = 0;
assign in27[17] = 0;
assign in27[18] = 0;
assign in27[19] = 0;
assign in27[20] = 0;
assign in27[21] = 0;
assign in27[22] = 0;
assign in27[23] = 0;
assign in27[24] = 0;
assign in27[25] = 0;
assign in27[26] = 0;
assign in28[31:28] = data_operandA[3:0];
assign in28[0] = 0;
assign in28[1] = 0;
assign in28[2] = 0;
assign in28[3] = 0;
assign in28[4] = 0;
assign in28[5] = 0;
assign in28[6] = 0;
assign in28[7] = 0;
assign in28[8] = 0;
assign in28[9] = 0;
assign in28[10] = 0;
assign in28[11] = 0;
assign in28[12] = 0;
assign in28[13] = 0;
assign in28[14] = 0;
assign in28[15] = 0;
assign in28[16] = 0;
assign in28[17] = 0;
assign in28[18] = 0;
assign in28[19] = 0;
assign in28[20] = 0;
assign in28[21] = 0;
assign in28[22] = 0;
assign in28[23] = 0;
assign in28[24] = 0;
assign in28[25] = 0;
assign in28[26] = 0;
assign in28[27] = 0;
assign in29[31:29] = data_operandA[2:0];
assign in29[0] = 0;
assign in29[1] = 0;
assign in29[2] = 0;
assign in29[3] = 0;
assign in29[4] = 0;
assign in29[5] = 0;
assign in29[6] = 0;
assign in29[7] = 0;
assign in29[8] = 0;
assign in29[9] = 0;
assign in29[10] = 0;
assign in29[11] = 0;
assign in29[12] = 0;
assign in29[13] = 0;
assign in29[14] = 0;
assign in29[15] = 0;
assign in29[16] = 0;
assign in29[17] = 0;
assign in29[18] = 0;
assign in29[19] = 0;
assign in29[20] = 0;
assign in29[21] = 0;
assign in29[22] = 0;
assign in29[23] = 0;
assign in29[24] = 0;
assign in29[25] = 0;
assign in29[26] = 0;
assign in29[27] = 0;
assign in29[28] = 0;
assign in30[31:30] = data_operandA[1:0];
assign in30[0] = 0;
assign in30[1] = 0;
assign in30[2] = 0;
assign in30[3] = 0;
assign in30[4] = 0;
assign in30[5] = 0;
assign in30[6] = 0;
assign in30[7] = 0;
assign in30[8] = 0;
assign in30[9] = 0;
assign in30[10] = 0;
assign in30[11] = 0;
assign in30[12] = 0;
assign in30[13] = 0;
assign in30[14] = 0;
assign in30[15] = 0;
assign in30[16] = 0;
assign in30[17] = 0;
assign in30[18] = 0;
assign in30[19] = 0;
assign in30[20] = 0;
assign in30[21] = 0;
assign in30[22] = 0;
assign in30[23] = 0;
assign in30[24] = 0;
assign in30[25] = 0;
assign in30[26] = 0;
assign in30[27] = 0;
assign in30[28] = 0;
assign in30[29] = 0;
assign in31[31:31] = data_operandA[0:0];
assign in31[0] = 0;
assign in31[1] = 0;
assign in31[2] = 0;
assign in31[3] = 0;
assign in31[4] = 0;
assign in31[5] = 0;
assign in31[6] = 0;
assign in31[7] = 0;
assign in31[8] = 0;
assign in31[9] = 0;
assign in31[10] = 0;
assign in31[11] = 0;
assign in31[12] = 0;
assign in31[13] = 0;
assign in31[14] = 0;
assign in31[15] = 0;
assign in31[16] = 0;
assign in31[17] = 0;
assign in31[18] = 0;
assign in31[19] = 0;
assign in31[20] = 0;
assign in31[21] = 0;
assign in31[22] = 0;
assign in31[23] = 0;
assign in31[24] = 0;
assign in31[25] = 0;
assign in31[26] = 0;
assign in31[27] = 0;
assign in31[28] = 0;
assign in31[29] = 0;
assign in31[30] = 0;
endmodule
	
