module or_32(data_operandA, data_operandB, or_enable, or_output);

	input [31:0] data_operandA, data_operandB;
	input or_enable;
	wire [31:0] ors;
	output [31:0] or_output;
	
	or or_0(ors[0], data_operandA[0], data_operandB[0]);
	or or_1(ors[1], data_operandA[1], data_operandB[1]);
	or or_2(ors[2], data_operandA[2], data_operandB[2]);
	or or_3(ors[3], data_operandA[3], data_operandB[3]);
	or or_4(ors[4], data_operandA[4], data_operandB[4]);
	or or_5(ors[5], data_operandA[5], data_operandB[5]);
	or or_6(ors[6], data_operandA[6], data_operandB[6]);
	or or_7(ors[7], data_operandA[7], data_operandB[7]);
	or or_8(ors[8], data_operandA[8], data_operandB[8]);
	or or_9(ors[9], data_operandA[9], data_operandB[9]);
	or or_10(ors[10], data_operandA[10], data_operandB[10]);
	or or_11(ors[11], data_operandA[11], data_operandB[11]);
	or or_12(ors[12], data_operandA[12], data_operandB[12]);
	or or_13(ors[13], data_operandA[13], data_operandB[13]);
	or or_14(ors[14], data_operandA[14], data_operandB[14]);
	or or_15(ors[15], data_operandA[15], data_operandB[15]);
	or or_16(ors[16], data_operandA[16], data_operandB[16]);
	or or_17(ors[17], data_operandA[17], data_operandB[17]);
	or or_18(ors[18], data_operandA[18], data_operandB[18]);
	or or_19(ors[19], data_operandA[19], data_operandB[19]);
	or or_20(ors[20], data_operandA[20], data_operandB[20]);
	or or_21(ors[21], data_operandA[21], data_operandB[21]);
	or or_22(ors[22], data_operandA[22], data_operandB[22]);
	or or_23(ors[23], data_operandA[23], data_operandB[23]);
	or or_24(ors[24], data_operandA[24], data_operandB[24]);
	or or_25(ors[25], data_operandA[25], data_operandB[25]);
	or or_26(ors[26], data_operandA[26], data_operandB[26]);
	or or_27(ors[27], data_operandA[27], data_operandB[27]);
	or or_28(ors[28], data_operandA[28], data_operandB[28]);
	or or_29(ors[29], data_operandA[29], data_operandB[29]);
	or or_30(ors[30], data_operandA[30], data_operandB[30]);
	or or_31(ors[31], data_operandA[31], data_operandB[31]);
	and and_0(or_output[0], ors[0], or_enable);
	and and_1(or_output[1], ors[1], or_enable);
	and and_2(or_output[2], ors[2], or_enable);
	and and_3(or_output[3], ors[3], or_enable);
	and and_4(or_output[4], ors[4], or_enable);
	and and_5(or_output[5], ors[5], or_enable);
	and and_6(or_output[6], ors[6], or_enable);
	and and_7(or_output[7], ors[7], or_enable);
	and and_8(or_output[8], ors[8], or_enable);
	and and_9(or_output[9], ors[9], or_enable);
	and and_10(or_output[10], ors[10], or_enable);
	and and_11(or_output[11], ors[11], or_enable);
	and and_12(or_output[12], ors[12], or_enable);
	and and_13(or_output[13], ors[13], or_enable);
	and and_14(or_output[14], ors[14], or_enable);
	and and_15(or_output[15], ors[15], or_enable);
	and and_16(or_output[16], ors[16], or_enable);
	and and_17(or_output[17], ors[17], or_enable);
	and and_18(or_output[18], ors[18], or_enable);
	and and_19(or_output[19], ors[19], or_enable);
	and and_20(or_output[20], ors[20], or_enable);
	and and_21(or_output[21], ors[21], or_enable);
	and and_22(or_output[22], ors[22], or_enable);
	and and_23(or_output[23], ors[23], or_enable);
	and and_24(or_output[24], ors[24], or_enable);
	and and_25(or_output[25], ors[25], or_enable);
	and and_26(or_output[26], ors[26], or_enable);
	and and_27(or_output[27], ors[27], or_enable);
	and and_28(or_output[28], ors[28], or_enable);
	and and_29(or_output[29], ors[29], or_enable);
	and and_30(or_output[30], ors[30], or_enable);
	and and_31(or_output[31], ors[31], or_enable);
	
endmodule
	