module tff16_tb;

endmodule