module cla(a, b, cin, g, p);

endmodule