module sra(data_operandA, ctrl_shiftamt, shifted_output, shift_enable);

	input [31:0] data_operandA;
	input [4:0] ctrl_shiftamt;
	input shift_enable;
	wire [31:0] muxed_output;
	output [31:0] shifted_output;
	
	
	wire [31:0] in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31;
	
	mux_32 mux_32_sra(muxed_output, ctrl_shiftamt, in0, in1, in2, in3, in4, in5, in6, in7, in8, in9, in10, in11, in12, in13, in14, in15, in16, in17, in18, in19, in20, in21, in22, in23, in24, in25, in26, in27, in28, in29, in30, in31);
	
	and and_0(shifted_output[0], muxed_output[0], shift_enable);
	and and_1(shifted_output[1], muxed_output[1], shift_enable);
	and and_2(shifted_output[2], muxed_output[2], shift_enable);
	and and_3(shifted_output[3], muxed_output[3], shift_enable);
	and and_4(shifted_output[4], muxed_output[4], shift_enable);
	and and_5(shifted_output[5], muxed_output[5], shift_enable);
	and and_6(shifted_output[6], muxed_output[6], shift_enable);
	and and_7(shifted_output[7], muxed_output[7], shift_enable);
	and and_8(shifted_output[8], muxed_output[8], shift_enable);
	and and_9(shifted_output[9], muxed_output[9], shift_enable);
	and and_10(shifted_output[10], muxed_output[10], shift_enable);
	and and_11(shifted_output[11], muxed_output[11], shift_enable);
	and and_12(shifted_output[12], muxed_output[12], shift_enable);
	and and_13(shifted_output[13], muxed_output[13], shift_enable);
	and and_14(shifted_output[14], muxed_output[14], shift_enable);
	and and_15(shifted_output[15], muxed_output[15], shift_enable);
	and and_16(shifted_output[16], muxed_output[16], shift_enable);
	and and_17(shifted_output[17], muxed_output[17], shift_enable);
	and and_18(shifted_output[18], muxed_output[18], shift_enable);
	and and_19(shifted_output[19], muxed_output[19], shift_enable);
	and and_20(shifted_output[20], muxed_output[20], shift_enable);
	and and_21(shifted_output[21], muxed_output[21], shift_enable);
	and and_22(shifted_output[22], muxed_output[22], shift_enable);
	and and_23(shifted_output[23], muxed_output[23], shift_enable);
	and and_24(shifted_output[24], muxed_output[24], shift_enable);
	and and_25(shifted_output[25], muxed_output[25], shift_enable);
	and and_26(shifted_output[26], muxed_output[26], shift_enable);
	and and_27(shifted_output[27], muxed_output[27], shift_enable);
	and and_28(shifted_output[28], muxed_output[28], shift_enable);
	and and_29(shifted_output[29], muxed_output[29], shift_enable);
	and and_30(shifted_output[30], muxed_output[30], shift_enable);
	and and_31(shifted_output[31], muxed_output[31], shift_enable);
	
	
	
assign in0[31:0] = data_operandA[31:0];
assign in1[30:0] = data_operandA[31:1];
assign in1[31] = data_operandA[31];
assign in2[29:0] = data_operandA[31:2];
assign in2[31] = data_operandA[31];
assign in2[30] = data_operandA[31];
assign in3[28:0] = data_operandA[31:3];
assign in3[31] = data_operandA[31];
assign in3[30] = data_operandA[31];
assign in3[29] = data_operandA[31];
assign in4[27:0] = data_operandA[31:4];
assign in4[31] = data_operandA[31];
assign in4[30] = data_operandA[31];
assign in4[29] = data_operandA[31];
assign in4[28] = data_operandA[31];
assign in5[26:0] = data_operandA[31:5];
assign in5[31] = data_operandA[31];
assign in5[30] = data_operandA[31];
assign in5[29] = data_operandA[31];
assign in5[28] = data_operandA[31];
assign in5[27] = data_operandA[31];
assign in6[25:0] = data_operandA[31:6];
assign in6[31] = data_operandA[31];
assign in6[30] = data_operandA[31];
assign in6[29] = data_operandA[31];
assign in6[28] = data_operandA[31];
assign in6[27] = data_operandA[31];
assign in6[26] = data_operandA[31];
assign in7[24:0] = data_operandA[31:7];
assign in7[31] = data_operandA[31];
assign in7[30] = data_operandA[31];
assign in7[29] = data_operandA[31];
assign in7[28] = data_operandA[31];
assign in7[27] = data_operandA[31];
assign in7[26] = data_operandA[31];
assign in7[25] = data_operandA[31];
assign in8[23:0] = data_operandA[31:8];
assign in8[31] = data_operandA[31];
assign in8[30] = data_operandA[31];
assign in8[29] = data_operandA[31];
assign in8[28] = data_operandA[31];
assign in8[27] = data_operandA[31];
assign in8[26] = data_operandA[31];
assign in8[25] = data_operandA[31];
assign in8[24] = data_operandA[31];
assign in9[22:0] = data_operandA[31:9];
assign in9[31] = data_operandA[31];
assign in9[30] = data_operandA[31];
assign in9[29] = data_operandA[31];
assign in9[28] = data_operandA[31];
assign in9[27] = data_operandA[31];
assign in9[26] = data_operandA[31];
assign in9[25] = data_operandA[31];
assign in9[24] = data_operandA[31];
assign in9[23] = data_operandA[31];
assign in10[21:0] = data_operandA[31:10];
assign in10[31] = data_operandA[31];
assign in10[30] = data_operandA[31];
assign in10[29] = data_operandA[31];
assign in10[28] = data_operandA[31];
assign in10[27] = data_operandA[31];
assign in10[26] = data_operandA[31];
assign in10[25] = data_operandA[31];
assign in10[24] = data_operandA[31];
assign in10[23] = data_operandA[31];
assign in10[22] = data_operandA[31];
assign in11[20:0] = data_operandA[31:11];
assign in11[31] = data_operandA[31];
assign in11[30] = data_operandA[31];
assign in11[29] = data_operandA[31];
assign in11[28] = data_operandA[31];
assign in11[27] = data_operandA[31];
assign in11[26] = data_operandA[31];
assign in11[25] = data_operandA[31];
assign in11[24] = data_operandA[31];
assign in11[23] = data_operandA[31];
assign in11[22] = data_operandA[31];
assign in11[21] = data_operandA[31];
assign in12[19:0] = data_operandA[31:12];
assign in12[31] = data_operandA[31];
assign in12[30] = data_operandA[31];
assign in12[29] = data_operandA[31];
assign in12[28] = data_operandA[31];
assign in12[27] = data_operandA[31];
assign in12[26] = data_operandA[31];
assign in12[25] = data_operandA[31];
assign in12[24] = data_operandA[31];
assign in12[23] = data_operandA[31];
assign in12[22] = data_operandA[31];
assign in12[21] = data_operandA[31];
assign in12[20] = data_operandA[31];
assign in13[18:0] = data_operandA[31:13];
assign in13[31] = data_operandA[31];
assign in13[30] = data_operandA[31];
assign in13[29] = data_operandA[31];
assign in13[28] = data_operandA[31];
assign in13[27] = data_operandA[31];
assign in13[26] = data_operandA[31];
assign in13[25] = data_operandA[31];
assign in13[24] = data_operandA[31];
assign in13[23] = data_operandA[31];
assign in13[22] = data_operandA[31];
assign in13[21] = data_operandA[31];
assign in13[20] = data_operandA[31];
assign in13[19] = data_operandA[31];
assign in14[17:0] = data_operandA[31:14];
assign in14[31] = data_operandA[31];
assign in14[30] = data_operandA[31];
assign in14[29] = data_operandA[31];
assign in14[28] = data_operandA[31];
assign in14[27] = data_operandA[31];
assign in14[26] = data_operandA[31];
assign in14[25] = data_operandA[31];
assign in14[24] = data_operandA[31];
assign in14[23] = data_operandA[31];
assign in14[22] = data_operandA[31];
assign in14[21] = data_operandA[31];
assign in14[20] = data_operandA[31];
assign in14[19] = data_operandA[31];
assign in14[18] = data_operandA[31];
assign in15[16:0] = data_operandA[31:15];
assign in15[31] = data_operandA[31];
assign in15[30] = data_operandA[31];
assign in15[29] = data_operandA[31];
assign in15[28] = data_operandA[31];
assign in15[27] = data_operandA[31];
assign in15[26] = data_operandA[31];
assign in15[25] = data_operandA[31];
assign in15[24] = data_operandA[31];
assign in15[23] = data_operandA[31];
assign in15[22] = data_operandA[31];
assign in15[21] = data_operandA[31];
assign in15[20] = data_operandA[31];
assign in15[19] = data_operandA[31];
assign in15[18] = data_operandA[31];
assign in15[17] = data_operandA[31];
assign in16[15:0] = data_operandA[31:16];
assign in16[31] = data_operandA[31];
assign in16[30] = data_operandA[31];
assign in16[29] = data_operandA[31];
assign in16[28] = data_operandA[31];
assign in16[27] = data_operandA[31];
assign in16[26] = data_operandA[31];
assign in16[25] = data_operandA[31];
assign in16[24] = data_operandA[31];
assign in16[23] = data_operandA[31];
assign in16[22] = data_operandA[31];
assign in16[21] = data_operandA[31];
assign in16[20] = data_operandA[31];
assign in16[19] = data_operandA[31];
assign in16[18] = data_operandA[31];
assign in16[17] = data_operandA[31];
assign in16[16] = data_operandA[31];
assign in17[14:0] = data_operandA[31:17];
assign in17[31] = data_operandA[31];
assign in17[30] = data_operandA[31];
assign in17[29] = data_operandA[31];
assign in17[28] = data_operandA[31];
assign in17[27] = data_operandA[31];
assign in17[26] = data_operandA[31];
assign in17[25] = data_operandA[31];
assign in17[24] = data_operandA[31];
assign in17[23] = data_operandA[31];
assign in17[22] = data_operandA[31];
assign in17[21] = data_operandA[31];
assign in17[20] = data_operandA[31];
assign in17[19] = data_operandA[31];
assign in17[18] = data_operandA[31];
assign in17[17] = data_operandA[31];
assign in17[16] = data_operandA[31];
assign in17[15] = data_operandA[31];
assign in18[13:0] = data_operandA[31:18];
assign in18[31] = data_operandA[31];
assign in18[30] = data_operandA[31];
assign in18[29] = data_operandA[31];
assign in18[28] = data_operandA[31];
assign in18[27] = data_operandA[31];
assign in18[26] = data_operandA[31];
assign in18[25] = data_operandA[31];
assign in18[24] = data_operandA[31];
assign in18[23] = data_operandA[31];
assign in18[22] = data_operandA[31];
assign in18[21] = data_operandA[31];
assign in18[20] = data_operandA[31];
assign in18[19] = data_operandA[31];
assign in18[18] = data_operandA[31];
assign in18[17] = data_operandA[31];
assign in18[16] = data_operandA[31];
assign in18[15] = data_operandA[31];
assign in18[14] = data_operandA[31];
assign in19[12:0] = data_operandA[31:19];
assign in19[31] = data_operandA[31];
assign in19[30] = data_operandA[31];
assign in19[29] = data_operandA[31];
assign in19[28] = data_operandA[31];
assign in19[27] = data_operandA[31];
assign in19[26] = data_operandA[31];
assign in19[25] = data_operandA[31];
assign in19[24] = data_operandA[31];
assign in19[23] = data_operandA[31];
assign in19[22] = data_operandA[31];
assign in19[21] = data_operandA[31];
assign in19[20] = data_operandA[31];
assign in19[19] = data_operandA[31];
assign in19[18] = data_operandA[31];
assign in19[17] = data_operandA[31];
assign in19[16] = data_operandA[31];
assign in19[15] = data_operandA[31];
assign in19[14] = data_operandA[31];
assign in19[13] = data_operandA[31];
assign in20[11:0] = data_operandA[31:20];
assign in20[31] = data_operandA[31];
assign in20[30] = data_operandA[31];
assign in20[29] = data_operandA[31];
assign in20[28] = data_operandA[31];
assign in20[27] = data_operandA[31];
assign in20[26] = data_operandA[31];
assign in20[25] = data_operandA[31];
assign in20[24] = data_operandA[31];
assign in20[23] = data_operandA[31];
assign in20[22] = data_operandA[31];
assign in20[21] = data_operandA[31];
assign in20[20] = data_operandA[31];
assign in20[19] = data_operandA[31];
assign in20[18] = data_operandA[31];
assign in20[17] = data_operandA[31];
assign in20[16] = data_operandA[31];
assign in20[15] = data_operandA[31];
assign in20[14] = data_operandA[31];
assign in20[13] = data_operandA[31];
assign in20[12] = data_operandA[31];
assign in21[10:0] = data_operandA[31:21];
assign in21[31] = data_operandA[31];
assign in21[30] = data_operandA[31];
assign in21[29] = data_operandA[31];
assign in21[28] = data_operandA[31];
assign in21[27] = data_operandA[31];
assign in21[26] = data_operandA[31];
assign in21[25] = data_operandA[31];
assign in21[24] = data_operandA[31];
assign in21[23] = data_operandA[31];
assign in21[22] = data_operandA[31];
assign in21[21] = data_operandA[31];
assign in21[20] = data_operandA[31];
assign in21[19] = data_operandA[31];
assign in21[18] = data_operandA[31];
assign in21[17] = data_operandA[31];
assign in21[16] = data_operandA[31];
assign in21[15] = data_operandA[31];
assign in21[14] = data_operandA[31];
assign in21[13] = data_operandA[31];
assign in21[12] = data_operandA[31];
assign in21[11] = data_operandA[31];
assign in22[9:0] = data_operandA[31:22];
assign in22[31] = data_operandA[31];
assign in22[30] = data_operandA[31];
assign in22[29] = data_operandA[31];
assign in22[28] = data_operandA[31];
assign in22[27] = data_operandA[31];
assign in22[26] = data_operandA[31];
assign in22[25] = data_operandA[31];
assign in22[24] = data_operandA[31];
assign in22[23] = data_operandA[31];
assign in22[22] = data_operandA[31];
assign in22[21] = data_operandA[31];
assign in22[20] = data_operandA[31];
assign in22[19] = data_operandA[31];
assign in22[18] = data_operandA[31];
assign in22[17] = data_operandA[31];
assign in22[16] = data_operandA[31];
assign in22[15] = data_operandA[31];
assign in22[14] = data_operandA[31];
assign in22[13] = data_operandA[31];
assign in22[12] = data_operandA[31];
assign in22[11] = data_operandA[31];
assign in22[10] = data_operandA[31];
assign in23[8:0] = data_operandA[31:23];
assign in23[31] = data_operandA[31];
assign in23[30] = data_operandA[31];
assign in23[29] = data_operandA[31];
assign in23[28] = data_operandA[31];
assign in23[27] = data_operandA[31];
assign in23[26] = data_operandA[31];
assign in23[25] = data_operandA[31];
assign in23[24] = data_operandA[31];
assign in23[23] = data_operandA[31];
assign in23[22] = data_operandA[31];
assign in23[21] = data_operandA[31];
assign in23[20] = data_operandA[31];
assign in23[19] = data_operandA[31];
assign in23[18] = data_operandA[31];
assign in23[17] = data_operandA[31];
assign in23[16] = data_operandA[31];
assign in23[15] = data_operandA[31];
assign in23[14] = data_operandA[31];
assign in23[13] = data_operandA[31];
assign in23[12] = data_operandA[31];
assign in23[11] = data_operandA[31];
assign in23[10] = data_operandA[31];
assign in23[9] = data_operandA[31];
assign in24[7:0] = data_operandA[31:24];
assign in24[31] = data_operandA[31];
assign in24[30] = data_operandA[31];
assign in24[29] = data_operandA[31];
assign in24[28] = data_operandA[31];
assign in24[27] = data_operandA[31];
assign in24[26] = data_operandA[31];
assign in24[25] = data_operandA[31];
assign in24[24] = data_operandA[31];
assign in24[23] = data_operandA[31];
assign in24[22] = data_operandA[31];
assign in24[21] = data_operandA[31];
assign in24[20] = data_operandA[31];
assign in24[19] = data_operandA[31];
assign in24[18] = data_operandA[31];
assign in24[17] = data_operandA[31];
assign in24[16] = data_operandA[31];
assign in24[15] = data_operandA[31];
assign in24[14] = data_operandA[31];
assign in24[13] = data_operandA[31];
assign in24[12] = data_operandA[31];
assign in24[11] = data_operandA[31];
assign in24[10] = data_operandA[31];
assign in24[9] = data_operandA[31];
assign in24[8] = data_operandA[31];
assign in25[6:0] = data_operandA[31:25];
assign in25[31] = data_operandA[31];
assign in25[30] = data_operandA[31];
assign in25[29] = data_operandA[31];
assign in25[28] = data_operandA[31];
assign in25[27] = data_operandA[31];
assign in25[26] = data_operandA[31];
assign in25[25] = data_operandA[31];
assign in25[24] = data_operandA[31];
assign in25[23] = data_operandA[31];
assign in25[22] = data_operandA[31];
assign in25[21] = data_operandA[31];
assign in25[20] = data_operandA[31];
assign in25[19] = data_operandA[31];
assign in25[18] = data_operandA[31];
assign in25[17] = data_operandA[31];
assign in25[16] = data_operandA[31];
assign in25[15] = data_operandA[31];
assign in25[14] = data_operandA[31];
assign in25[13] = data_operandA[31];
assign in25[12] = data_operandA[31];
assign in25[11] = data_operandA[31];
assign in25[10] = data_operandA[31];
assign in25[9] = data_operandA[31];
assign in25[8] = data_operandA[31];
assign in25[7] = data_operandA[31];
assign in26[5:0] = data_operandA[31:26];
assign in26[31] = data_operandA[31];
assign in26[30] = data_operandA[31];
assign in26[29] = data_operandA[31];
assign in26[28] = data_operandA[31];
assign in26[27] = data_operandA[31];
assign in26[26] = data_operandA[31];
assign in26[25] = data_operandA[31];
assign in26[24] = data_operandA[31];
assign in26[23] = data_operandA[31];
assign in26[22] = data_operandA[31];
assign in26[21] = data_operandA[31];
assign in26[20] = data_operandA[31];
assign in26[19] = data_operandA[31];
assign in26[18] = data_operandA[31];
assign in26[17] = data_operandA[31];
assign in26[16] = data_operandA[31];
assign in26[15] = data_operandA[31];
assign in26[14] = data_operandA[31];
assign in26[13] = data_operandA[31];
assign in26[12] = data_operandA[31];
assign in26[11] = data_operandA[31];
assign in26[10] = data_operandA[31];
assign in26[9] = data_operandA[31];
assign in26[8] = data_operandA[31];
assign in26[7] = data_operandA[31];
assign in26[6] = data_operandA[31];
assign in27[4:0] = data_operandA[31:27];
assign in27[31] = data_operandA[31];
assign in27[30] = data_operandA[31];
assign in27[29] = data_operandA[31];
assign in27[28] = data_operandA[31];
assign in27[27] = data_operandA[31];
assign in27[26] = data_operandA[31];
assign in27[25] = data_operandA[31];
assign in27[24] = data_operandA[31];
assign in27[23] = data_operandA[31];
assign in27[22] = data_operandA[31];
assign in27[21] = data_operandA[31];
assign in27[20] = data_operandA[31];
assign in27[19] = data_operandA[31];
assign in27[18] = data_operandA[31];
assign in27[17] = data_operandA[31];
assign in27[16] = data_operandA[31];
assign in27[15] = data_operandA[31];
assign in27[14] = data_operandA[31];
assign in27[13] = data_operandA[31];
assign in27[12] = data_operandA[31];
assign in27[11] = data_operandA[31];
assign in27[10] = data_operandA[31];
assign in27[9] = data_operandA[31];
assign in27[8] = data_operandA[31];
assign in27[7] = data_operandA[31];
assign in27[6] = data_operandA[31];
assign in27[5] = data_operandA[31];
assign in28[3:0] = data_operandA[31:28];
assign in28[31] = data_operandA[31];
assign in28[30] = data_operandA[31];
assign in28[29] = data_operandA[31];
assign in28[28] = data_operandA[31];
assign in28[27] = data_operandA[31];
assign in28[26] = data_operandA[31];
assign in28[25] = data_operandA[31];
assign in28[24] = data_operandA[31];
assign in28[23] = data_operandA[31];
assign in28[22] = data_operandA[31];
assign in28[21] = data_operandA[31];
assign in28[20] = data_operandA[31];
assign in28[19] = data_operandA[31];
assign in28[18] = data_operandA[31];
assign in28[17] = data_operandA[31];
assign in28[16] = data_operandA[31];
assign in28[15] = data_operandA[31];
assign in28[14] = data_operandA[31];
assign in28[13] = data_operandA[31];
assign in28[12] = data_operandA[31];
assign in28[11] = data_operandA[31];
assign in28[10] = data_operandA[31];
assign in28[9] = data_operandA[31];
assign in28[8] = data_operandA[31];
assign in28[7] = data_operandA[31];
assign in28[6] = data_operandA[31];
assign in28[5] = data_operandA[31];
assign in28[4] = data_operandA[31];
assign in29[2:0] = data_operandA[31:29];
assign in29[31] = data_operandA[31];
assign in29[30] = data_operandA[31];
assign in29[29] = data_operandA[31];
assign in29[28] = data_operandA[31];
assign in29[27] = data_operandA[31];
assign in29[26] = data_operandA[31];
assign in29[25] = data_operandA[31];
assign in29[24] = data_operandA[31];
assign in29[23] = data_operandA[31];
assign in29[22] = data_operandA[31];
assign in29[21] = data_operandA[31];
assign in29[20] = data_operandA[31];
assign in29[19] = data_operandA[31];
assign in29[18] = data_operandA[31];
assign in29[17] = data_operandA[31];
assign in29[16] = data_operandA[31];
assign in29[15] = data_operandA[31];
assign in29[14] = data_operandA[31];
assign in29[13] = data_operandA[31];
assign in29[12] = data_operandA[31];
assign in29[11] = data_operandA[31];
assign in29[10] = data_operandA[31];
assign in29[9] = data_operandA[31];
assign in29[8] = data_operandA[31];
assign in29[7] = data_operandA[31];
assign in29[6] = data_operandA[31];
assign in29[5] = data_operandA[31];
assign in29[4] = data_operandA[31];
assign in29[3] = data_operandA[31];
assign in30[1:0] = data_operandA[31:30];
assign in30[31] = data_operandA[31];
assign in30[30] = data_operandA[31];
assign in30[29] = data_operandA[31];
assign in30[28] = data_operandA[31];
assign in30[27] = data_operandA[31];
assign in30[26] = data_operandA[31];
assign in30[25] = data_operandA[31];
assign in30[24] = data_operandA[31];
assign in30[23] = data_operandA[31];
assign in30[22] = data_operandA[31];
assign in30[21] = data_operandA[31];
assign in30[20] = data_operandA[31];
assign in30[19] = data_operandA[31];
assign in30[18] = data_operandA[31];
assign in30[17] = data_operandA[31];
assign in30[16] = data_operandA[31];
assign in30[15] = data_operandA[31];
assign in30[14] = data_operandA[31];
assign in30[13] = data_operandA[31];
assign in30[12] = data_operandA[31];
assign in30[11] = data_operandA[31];
assign in30[10] = data_operandA[31];
assign in30[9] = data_operandA[31];
assign in30[8] = data_operandA[31];
assign in30[7] = data_operandA[31];
assign in30[6] = data_operandA[31];
assign in30[5] = data_operandA[31];
assign in30[4] = data_operandA[31];
assign in30[3] = data_operandA[31];
assign in30[2] = data_operandA[31];
assign in31[0:0] = data_operandA[31:31];
assign in31[31] = data_operandA[31];
assign in31[30] = data_operandA[31];
assign in31[29] = data_operandA[31];
assign in31[28] = data_operandA[31];
assign in31[27] = data_operandA[31];
assign in31[26] = data_operandA[31];
assign in31[25] = data_operandA[31];
assign in31[24] = data_operandA[31];
assign in31[23] = data_operandA[31];
assign in31[22] = data_operandA[31];
assign in31[21] = data_operandA[31];
assign in31[20] = data_operandA[31];
assign in31[19] = data_operandA[31];
assign in31[18] = data_operandA[31];
assign in31[17] = data_operandA[31];
assign in31[16] = data_operandA[31];
assign in31[15] = data_operandA[31];
assign in31[14] = data_operandA[31];
assign in31[13] = data_operandA[31];
assign in31[12] = data_operandA[31];
assign in31[11] = data_operandA[31];
assign in31[10] = data_operandA[31];
assign in31[9] = data_operandA[31];
assign in31[8] = data_operandA[31];
assign in31[7] = data_operandA[31];
assign in31[6] = data_operandA[31];
assign in31[5] = data_operandA[31];
assign in31[4] = data_operandA[31];
assign in31[3] = data_operandA[31];
assign in31[2] = data_operandA[31];
assign in31[1] = data_operandA[31];
	
endmodule