module less_than(A, B, out);

	input [31:0] A, B;
	output out;
	
	

endmodule