module not_32(A, Out);

	input [31:0] A;
	output [31:0] Out;
	
	not not0(Out[0], A[0]);
	not not1(Out[1], A[1]);
	not not2(Out[2], A[2]);
	not not3(Out[3], A[3]);
	not not4(Out[4], A[4]);
	not not5(Out[5], A[5]);
	not not6(Out[6], A[6]);
	not not7(Out[7], A[7]);
	not not8(Out[8], A[8]);
	not not9(Out[9], A[9]);
	not not10(Out[10], A[10]);
	not not11(Out[11], A[11]);
	not not12(Out[12], A[12]);
	not not13(Out[13], A[13]);
	not not14(Out[14], A[14]);
	not not15(Out[15], A[15]);
	not not16(Out[16], A[16]);
	not not17(Out[17], A[17]);
	not not18(Out[18], A[18]);
	not not19(Out[19], A[19]);
	not not20(Out[20], A[20]);
	not not21(Out[21], A[21]);
	not not22(Out[22], A[22]);
	not not23(Out[23], A[23]);
	not not24(Out[24], A[24]);
	not not25(Out[25], A[25]);
	not not26(Out[26], A[26]);
	not not27(Out[27], A[27]);
	not not28(Out[28], A[28]);
	not not29(Out[29], A[29]);
	not not30(Out[30], A[30]);
	not not31(Out[31], A[31]);

endmodule